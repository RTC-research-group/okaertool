
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package okt_top_pkg is
	constant ROME_DATA_BITS_WIDTH      : integer := 8;
	constant NODE_DATA_BITS_WIDTH      : integer := 8;
	constant SPINNAKER_BITS_DATA_WIDTH : integer := 8;
	constant COMMAND_BIT_WIDTH         : integer := 5;
	constant OUT_DATA_BITS_WIDTH       : integer := 16;
	constant CONFIG_BITS_WIDTH         : integer := 16;
	constant CONFIG_NUN_DEVICES        : integer := 2;

end okt_top_pkg;

package body okt_top_pkg is

end okt_top_pkg;
